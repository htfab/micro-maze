`default_nettype none

module maze_data (
    input wire [3:0] x,
    input wire [3:0] x_alt,
    input wire [3:0] y,
    input wire [3:0] y_alt,
    output reg horizontal,
    output reg vertical
);

always @(*) begin
    case({y_alt, x})
        8'b0000_0000: horizontal = 1'b1;
        8'b0000_0001: horizontal = 1'b1;
        8'b0000_0010: horizontal = 1'b1;
        8'b0000_0011: horizontal = 1'b1;
        8'b0000_0100: horizontal = 1'b1;
        8'b0000_0101: horizontal = 1'b1;
        8'b0000_0110: horizontal = 1'b1;
        8'b0000_0111: horizontal = 1'b1;
        8'b0000_1000: horizontal = 1'b1;
        8'b0000_1001: horizontal = 1'b1;
        8'b0000_1010: horizontal = 1'bx;
        8'b0000_1011: horizontal = 1'bx;
        8'b0000_1100: horizontal = 1'bx;
        8'b0000_1101: horizontal = 1'bx;
        8'b0000_1110: horizontal = 1'bx;
        8'b0000_1111: horizontal = 1'bx;

        8'b0001_0000: horizontal = 1'b0;
        8'b0001_0001: horizontal = 1'b1;
        8'b0001_0010: horizontal = 1'b1;
        8'b0001_0011: horizontal = 1'b0;
        8'b0001_0100: horizontal = 1'b0;
        8'b0001_0101: horizontal = 1'b0;
        8'b0001_0110: horizontal = 1'b1;
        8'b0001_0111: horizontal = 1'b1;
        8'b0001_1000: horizontal = 1'b0;
        8'b0001_1001: horizontal = 1'b0;
        8'b0001_1010: horizontal = 1'bx;
        8'b0001_1011: horizontal = 1'bx;
        8'b0001_1100: horizontal = 1'bx;
        8'b0001_1101: horizontal = 1'bx;
        8'b0001_1110: horizontal = 1'bx;
        8'b0001_1111: horizontal = 1'bx;

        8'b0010_0000: horizontal = 1'b0;
        8'b0010_0001: horizontal = 1'b1;
        8'b0010_0010: horizontal = 1'b0;
        8'b0010_0011: horizontal = 1'b1;
        8'b0010_0100: horizontal = 1'b0;
        8'b0010_0101: horizontal = 1'b0;
        8'b0010_0110: horizontal = 1'b0;
        8'b0010_0111: horizontal = 1'b1;
        8'b0010_1000: horizontal = 1'b1;
        8'b0010_1001: horizontal = 1'b0;
        8'b0010_1010: horizontal = 1'bx;
        8'b0010_1011: horizontal = 1'bx;
        8'b0010_1100: horizontal = 1'bx;
        8'b0010_1101: horizontal = 1'bx;
        8'b0010_1110: horizontal = 1'bx;
        8'b0010_1111: horizontal = 1'bx;

        8'b0011_0000: horizontal = 1'b0;
        8'b0011_0001: horizontal = 1'b0;
        8'b0011_0010: horizontal = 1'b1;
        8'b0011_0011: horizontal = 1'b1;
        8'b0011_0100: horizontal = 1'b1;
        8'b0011_0101: horizontal = 1'b0;
        8'b0011_0110: horizontal = 1'b0;
        8'b0011_0111: horizontal = 1'b0;
        8'b0011_1000: horizontal = 1'b0;
        8'b0011_1001: horizontal = 1'b0;
        8'b0011_1010: horizontal = 1'bx;
        8'b0011_1011: horizontal = 1'bx;
        8'b0011_1100: horizontal = 1'bx;
        8'b0011_1101: horizontal = 1'bx;
        8'b0011_1110: horizontal = 1'bx;
        8'b0011_1111: horizontal = 1'bx;

        8'b0100_0000: horizontal = 1'b0;
        8'b0100_0001: horizontal = 1'b0;
        8'b0100_0010: horizontal = 1'b1;
        8'b0100_0011: horizontal = 1'b1;
        8'b0100_0100: horizontal = 1'b0;
        8'b0100_0101: horizontal = 1'b0;
        8'b0100_0110: horizontal = 1'b1;
        8'b0100_0111: horizontal = 1'b1;
        8'b0100_1000: horizontal = 1'b1;
        8'b0100_1001: horizontal = 1'b1;
        8'b0100_1010: horizontal = 1'bx;
        8'b0100_1011: horizontal = 1'bx;
        8'b0100_1100: horizontal = 1'bx;
        8'b0100_1101: horizontal = 1'bx;
        8'b0100_1110: horizontal = 1'bx;
        8'b0100_1111: horizontal = 1'bx;

        8'b0101_0000: horizontal = 1'b1;
        8'b0101_0001: horizontal = 1'b1;
        8'b0101_0010: horizontal = 1'b0;
        8'b0101_0011: horizontal = 1'b1;
        8'b0101_0100: horizontal = 1'b1;
        8'b0101_0101: horizontal = 1'b1;
        8'b0101_0110: horizontal = 1'b1;
        8'b0101_0111: horizontal = 1'b1;
        8'b0101_1000: horizontal = 1'b1;
        8'b0101_1001: horizontal = 1'b1;
        8'b0101_1010: horizontal = 1'bx;
        8'b0101_1011: horizontal = 1'bx;
        8'b0101_1100: horizontal = 1'bx;
        8'b0101_1101: horizontal = 1'bx;
        8'b0101_1110: horizontal = 1'bx;
        8'b0101_1111: horizontal = 1'bx;

        8'b0110_0000: horizontal = 1'b0;
        8'b0110_0001: horizontal = 1'b0;
        8'b0110_0010: horizontal = 1'b1;
        8'b0110_0011: horizontal = 1'b0;
        8'b0110_0100: horizontal = 1'b0;
        8'b0110_0101: horizontal = 1'b0;
        8'b0110_0110: horizontal = 1'b0;
        8'b0110_0111: horizontal = 1'b1;
        8'b0110_1000: horizontal = 1'b1;
        8'b0110_1001: horizontal = 1'b0;
        8'b0110_1010: horizontal = 1'bx;
        8'b0110_1011: horizontal = 1'bx;
        8'b0110_1100: horizontal = 1'bx;
        8'b0110_1101: horizontal = 1'bx;
        8'b0110_1110: horizontal = 1'bx;
        8'b0110_1111: horizontal = 1'bx;

        8'b0111_0000: horizontal = 1'b0;
        8'b0111_0001: horizontal = 1'b1;
        8'b0111_0010: horizontal = 1'b1;
        8'b0111_0011: horizontal = 1'b0;
        8'b0111_0100: horizontal = 1'b0;
        8'b0111_0101: horizontal = 1'b0;
        8'b0111_0110: horizontal = 1'b0;
        8'b0111_0111: horizontal = 1'b1;
        8'b0111_1000: horizontal = 1'b1;
        8'b0111_1001: horizontal = 1'b0;
        8'b0111_1010: horizontal = 1'bx;
        8'b0111_1011: horizontal = 1'bx;
        8'b0111_1100: horizontal = 1'bx;
        8'b0111_1101: horizontal = 1'bx;
        8'b0111_1110: horizontal = 1'bx;
        8'b0111_1111: horizontal = 1'bx;

        8'b1000_0000: horizontal = 1'b0;
        8'b1000_0001: horizontal = 1'b0;
        8'b1000_0010: horizontal = 1'b1;
        8'b1000_0011: horizontal = 1'b1;
        8'b1000_0100: horizontal = 1'b1;
        8'b1000_0101: horizontal = 1'b1;
        8'b1000_0110: horizontal = 1'b1;
        8'b1000_0111: horizontal = 1'b0;
        8'b1000_1000: horizontal = 1'b0;
        8'b1000_1001: horizontal = 1'b0;
        8'b1000_1010: horizontal = 1'bx;
        8'b1000_1011: horizontal = 1'bx;
        8'b1000_1100: horizontal = 1'bx;
        8'b1000_1101: horizontal = 1'bx;
        8'b1000_1110: horizontal = 1'bx;
        8'b1000_1111: horizontal = 1'bx;

        8'b1001_0000: horizontal = 1'b0;
        8'b1001_0001: horizontal = 1'b0;
        8'b1001_0010: horizontal = 1'b1;
        8'b1001_0011: horizontal = 1'b1;
        8'b1001_0100: horizontal = 1'b0;
        8'b1001_0101: horizontal = 1'b1;
        8'b1001_0110: horizontal = 1'b1;
        8'b1001_0111: horizontal = 1'b1;
        8'b1001_1000: horizontal = 1'b0;
        8'b1001_1001: horizontal = 1'b0;
        8'b1001_1010: horizontal = 1'bx;
        8'b1001_1011: horizontal = 1'bx;
        8'b1001_1100: horizontal = 1'bx;
        8'b1001_1101: horizontal = 1'bx;
        8'b1001_1110: horizontal = 1'bx;
        8'b1001_1111: horizontal = 1'bx;

        8'b1010_0000: horizontal = 1'b1;
        8'b1010_0001: horizontal = 1'b1;
        8'b1010_0010: horizontal = 1'b1;
        8'b1010_0011: horizontal = 1'b1;
        8'b1010_0100: horizontal = 1'b1;
        8'b1010_0101: horizontal = 1'b1;
        8'b1010_0110: horizontal = 1'b1;
        8'b1010_0111: horizontal = 1'b1;
        8'b1010_1000: horizontal = 1'b1;
        8'b1010_1001: horizontal = 1'b1;
        8'b1010_1010: horizontal = 1'bx;
        8'b1010_1011: horizontal = 1'bx;
        8'b1010_1100: horizontal = 1'bx;
        8'b1010_1101: horizontal = 1'bx;
        8'b1010_1110: horizontal = 1'bx;
        8'b1010_1111: horizontal = 1'bx;

        8'b1011_0000: horizontal = 1'bx;
        8'b1011_0001: horizontal = 1'bx;
        8'b1011_0010: horizontal = 1'bx;
        8'b1011_0011: horizontal = 1'bx;
        8'b1011_0100: horizontal = 1'bx;
        8'b1011_0101: horizontal = 1'bx;
        8'b1011_0110: horizontal = 1'bx;
        8'b1011_0111: horizontal = 1'bx;
        8'b1011_1000: horizontal = 1'bx;
        8'b1011_1001: horizontal = 1'bx;
        8'b1011_1010: horizontal = 1'bx;
        8'b1011_1011: horizontal = 1'bx;
        8'b1011_1100: horizontal = 1'bx;
        8'b1011_1101: horizontal = 1'bx;
        8'b1011_1110: horizontal = 1'bx;
        8'b1011_1111: horizontal = 1'bx;

        8'b1100_0000: horizontal = 1'bx;
        8'b1100_0001: horizontal = 1'bx;
        8'b1100_0010: horizontal = 1'bx;
        8'b1100_0011: horizontal = 1'bx;
        8'b1100_0100: horizontal = 1'bx;
        8'b1100_0101: horizontal = 1'bx;
        8'b1100_0110: horizontal = 1'bx;
        8'b1100_0111: horizontal = 1'bx;
        8'b1100_1000: horizontal = 1'bx;
        8'b1100_1001: horizontal = 1'bx;
        8'b1100_1010: horizontal = 1'bx;
        8'b1100_1011: horizontal = 1'bx;
        8'b1100_1100: horizontal = 1'bx;
        8'b1100_1101: horizontal = 1'bx;
        8'b1100_1110: horizontal = 1'bx;
        8'b1100_1111: horizontal = 1'bx;

        8'b1101_0000: horizontal = 1'bx;
        8'b1101_0001: horizontal = 1'bx;
        8'b1101_0010: horizontal = 1'bx;
        8'b1101_0011: horizontal = 1'bx;
        8'b1101_0100: horizontal = 1'bx;
        8'b1101_0101: horizontal = 1'bx;
        8'b1101_0110: horizontal = 1'bx;
        8'b1101_0111: horizontal = 1'bx;
        8'b1101_1000: horizontal = 1'bx;
        8'b1101_1001: horizontal = 1'bx;
        8'b1101_1010: horizontal = 1'bx;
        8'b1101_1011: horizontal = 1'bx;
        8'b1101_1100: horizontal = 1'bx;
        8'b1101_1101: horizontal = 1'bx;
        8'b1101_1110: horizontal = 1'bx;
        8'b1101_1111: horizontal = 1'bx;

        8'b1110_0000: horizontal = 1'bx;
        8'b1110_0001: horizontal = 1'bx;
        8'b1110_0010: horizontal = 1'bx;
        8'b1110_0011: horizontal = 1'bx;
        8'b1110_0100: horizontal = 1'bx;
        8'b1110_0101: horizontal = 1'bx;
        8'b1110_0110: horizontal = 1'bx;
        8'b1110_0111: horizontal = 1'bx;
        8'b1110_1000: horizontal = 1'bx;
        8'b1110_1001: horizontal = 1'bx;
        8'b1110_1010: horizontal = 1'bx;
        8'b1110_1011: horizontal = 1'bx;
        8'b1110_1100: horizontal = 1'bx;
        8'b1110_1101: horizontal = 1'bx;
        8'b1110_1110: horizontal = 1'bx;
        8'b1110_1111: horizontal = 1'bx;

        8'b1111_0000: horizontal = 1'bx;
        8'b1111_0001: horizontal = 1'bx;
        8'b1111_0010: horizontal = 1'bx;
        8'b1111_0011: horizontal = 1'bx;
        8'b1111_0100: horizontal = 1'bx;
        8'b1111_0101: horizontal = 1'bx;
        8'b1111_0110: horizontal = 1'bx;
        8'b1111_0111: horizontal = 1'bx;
        8'b1111_1000: horizontal = 1'bx;
        8'b1111_1001: horizontal = 1'bx;
        8'b1111_1010: horizontal = 1'bx;
        8'b1111_1011: horizontal = 1'bx;
        8'b1111_1100: horizontal = 1'bx;
        8'b1111_1101: horizontal = 1'bx;
        8'b1111_1110: horizontal = 1'bx;
        8'b1111_1111: horizontal = 1'bx;

    endcase
    case({y, x_alt})
        8'b0000_0000: vertical = 1'b1;
        8'b0000_0001: vertical = 1'b0;
        8'b0000_0010: vertical = 1'b0;
        8'b0000_0011: vertical = 1'b0;
        8'b0000_0100: vertical = 1'b1;
        8'b0000_0101: vertical = 1'b0;
        8'b0000_0110: vertical = 1'b0;
        8'b0000_0111: vertical = 1'b0;
        8'b0000_1000: vertical = 1'b0;
        8'b0000_1001: vertical = 1'b1;
        8'b0000_1010: vertical = 1'b1;
        8'b0000_1011: vertical = 1'bx;
        8'b0000_1100: vertical = 1'bx;
        8'b0000_1101: vertical = 1'bx;
        8'b0000_1110: vertical = 1'bx;
        8'b0000_1111: vertical = 1'bx;

        8'b0001_0000: vertical = 1'b1;
        8'b0001_0001: vertical = 1'b0;
        8'b0001_0010: vertical = 1'b0;
        8'b0001_0011: vertical = 1'b1;
        8'b0001_0100: vertical = 1'b1;
        8'b0001_0101: vertical = 1'b1;
        8'b0001_0110: vertical = 1'b1;
        8'b0001_0111: vertical = 1'b0;
        8'b0001_1000: vertical = 1'b1;
        8'b0001_1001: vertical = 1'b0;
        8'b0001_1010: vertical = 1'b1;
        8'b0001_1011: vertical = 1'bx;
        8'b0001_1100: vertical = 1'bx;
        8'b0001_1101: vertical = 1'bx;
        8'b0001_1110: vertical = 1'bx;
        8'b0001_1111: vertical = 1'bx;

        8'b0010_0000: vertical = 1'b1;
        8'b0010_0001: vertical = 1'b1;
        8'b0010_0010: vertical = 1'b1;
        8'b0010_0011: vertical = 1'b0;
        8'b0010_0100: vertical = 1'b0;
        8'b0010_0101: vertical = 1'b1;
        8'b0010_0110: vertical = 1'b1;
        8'b0010_0111: vertical = 1'b1;
        8'b0010_1000: vertical = 1'b0;
        8'b0010_1001: vertical = 1'b1;
        8'b0010_1010: vertical = 1'b1;
        8'b0010_1011: vertical = 1'bx;
        8'b0010_1100: vertical = 1'bx;
        8'b0010_1101: vertical = 1'bx;
        8'b0010_1110: vertical = 1'bx;
        8'b0010_1111: vertical = 1'bx;

        8'b0011_0000: vertical = 1'b1;
        8'b0011_0001: vertical = 1'b1;
        8'b0011_0010: vertical = 1'b0;
        8'b0011_0011: vertical = 1'b0;
        8'b0011_0100: vertical = 1'b0;
        8'b0011_0101: vertical = 1'b1;
        8'b0011_0110: vertical = 1'b1;
        8'b0011_0111: vertical = 1'b0;
        8'b0011_1000: vertical = 1'b1;
        8'b0011_1001: vertical = 1'b0;
        8'b0011_1010: vertical = 1'b1;
        8'b0011_1011: vertical = 1'bx;
        8'b0011_1100: vertical = 1'bx;
        8'b0011_1101: vertical = 1'bx;
        8'b0011_1110: vertical = 1'bx;
        8'b0011_1111: vertical = 1'bx;

        8'b0100_0000: vertical = 1'b1;
        8'b0100_0001: vertical = 1'b0;
        8'b0100_0010: vertical = 1'b1;
        8'b0100_0011: vertical = 1'b0;
        8'b0100_0100: vertical = 1'b0;
        8'b0100_0101: vertical = 1'b1;
        8'b0100_0110: vertical = 1'b0;
        8'b0100_0111: vertical = 1'b0;
        8'b0100_1000: vertical = 1'b0;
        8'b0100_1001: vertical = 1'b0;
        8'b0100_1010: vertical = 1'b1;
        8'b0100_1011: vertical = 1'bx;
        8'b0100_1100: vertical = 1'bx;
        8'b0100_1101: vertical = 1'bx;
        8'b0100_1110: vertical = 1'bx;
        8'b0100_1111: vertical = 1'bx;

        8'b0101_0000: vertical = 1'b1;
        8'b0101_0001: vertical = 1'b0;
        8'b0101_0010: vertical = 1'b1;
        8'b0101_0011: vertical = 1'b0;
        8'b0101_0100: vertical = 1'b1;
        8'b0101_0101: vertical = 1'b0;
        8'b0101_0110: vertical = 1'b1;
        8'b0101_0111: vertical = 1'b0;
        8'b0101_1000: vertical = 1'b0;
        8'b0101_1001: vertical = 1'b0;
        8'b0101_1010: vertical = 1'b1;
        8'b0101_1011: vertical = 1'bx;
        8'b0101_1100: vertical = 1'bx;
        8'b0101_1101: vertical = 1'bx;
        8'b0101_1110: vertical = 1'bx;
        8'b0101_1111: vertical = 1'bx;

        8'b0110_0000: vertical = 1'b1;
        8'b0110_0001: vertical = 1'b1;
        8'b0110_0010: vertical = 1'b0;
        8'b0110_0011: vertical = 1'b1;
        8'b0110_0100: vertical = 1'b1;
        8'b0110_0101: vertical = 1'b1;
        8'b0110_0110: vertical = 1'b1;
        8'b0110_0111: vertical = 1'b0;
        8'b0110_1000: vertical = 1'b0;
        8'b0110_1001: vertical = 1'b1;
        8'b0110_1010: vertical = 1'b1;
        8'b0110_1011: vertical = 1'bx;
        8'b0110_1100: vertical = 1'bx;
        8'b0110_1101: vertical = 1'bx;
        8'b0110_1110: vertical = 1'bx;
        8'b0110_1111: vertical = 1'bx;

        8'b0111_0000: vertical = 1'b1;
        8'b0111_0001: vertical = 1'b1;
        8'b0111_0010: vertical = 1'b0;
        8'b0111_0011: vertical = 1'b0;
        8'b0111_0100: vertical = 1'b1;
        8'b0111_0101: vertical = 1'b1;
        8'b0111_0110: vertical = 1'b0;
        8'b0111_0111: vertical = 1'b0;
        8'b0111_1000: vertical = 1'b0;
        8'b0111_1001: vertical = 1'b1;
        8'b0111_1010: vertical = 1'b1;
        8'b0111_1011: vertical = 1'bx;
        8'b0111_1100: vertical = 1'bx;
        8'b0111_1101: vertical = 1'bx;
        8'b0111_1110: vertical = 1'bx;
        8'b0111_1111: vertical = 1'bx;

        8'b1000_0000: vertical = 1'b1;
        8'b1000_0001: vertical = 1'b1;
        8'b1000_0010: vertical = 1'b1;
        8'b1000_0011: vertical = 1'b0;
        8'b1000_0100: vertical = 1'b0;
        8'b1000_0101: vertical = 1'b0;
        8'b1000_0110: vertical = 1'b0;
        8'b1000_0111: vertical = 1'b0;
        8'b1000_1000: vertical = 1'b1;
        8'b1000_1001: vertical = 1'b1;
        8'b1000_1010: vertical = 1'b1;
        8'b1000_1011: vertical = 1'bx;
        8'b1000_1100: vertical = 1'bx;
        8'b1000_1101: vertical = 1'bx;
        8'b1000_1110: vertical = 1'bx;
        8'b1000_1111: vertical = 1'bx;

        8'b1001_0000: vertical = 1'b1;
        8'b1001_0001: vertical = 1'b0;
        8'b1001_0010: vertical = 1'b0;
        8'b1001_0011: vertical = 1'b0;
        8'b1001_0100: vertical = 1'b0;
        8'b1001_0101: vertical = 1'b1;
        8'b1001_0110: vertical = 1'b0;
        8'b1001_0111: vertical = 1'b0;
        8'b1001_1000: vertical = 1'b0;
        8'b1001_1001: vertical = 1'b1;
        8'b1001_1010: vertical = 1'b1;
        8'b1001_1011: vertical = 1'bx;
        8'b1001_1100: vertical = 1'bx;
        8'b1001_1101: vertical = 1'bx;
        8'b1001_1110: vertical = 1'bx;
        8'b1001_1111: vertical = 1'bx;

        8'b1010_0000: vertical = 1'bx;
        8'b1010_0001: vertical = 1'bx;
        8'b1010_0010: vertical = 1'bx;
        8'b1010_0011: vertical = 1'bx;
        8'b1010_0100: vertical = 1'bx;
        8'b1010_0101: vertical = 1'bx;
        8'b1010_0110: vertical = 1'bx;
        8'b1010_0111: vertical = 1'bx;
        8'b1010_1000: vertical = 1'bx;
        8'b1010_1001: vertical = 1'bx;
        8'b1010_1010: vertical = 1'bx;
        8'b1010_1011: vertical = 1'bx;
        8'b1010_1100: vertical = 1'bx;
        8'b1010_1101: vertical = 1'bx;
        8'b1010_1110: vertical = 1'bx;
        8'b1010_1111: vertical = 1'bx;

        8'b1011_0000: vertical = 1'bx;
        8'b1011_0001: vertical = 1'bx;
        8'b1011_0010: vertical = 1'bx;
        8'b1011_0011: vertical = 1'bx;
        8'b1011_0100: vertical = 1'bx;
        8'b1011_0101: vertical = 1'bx;
        8'b1011_0110: vertical = 1'bx;
        8'b1011_0111: vertical = 1'bx;
        8'b1011_1000: vertical = 1'bx;
        8'b1011_1001: vertical = 1'bx;
        8'b1011_1010: vertical = 1'bx;
        8'b1011_1011: vertical = 1'bx;
        8'b1011_1100: vertical = 1'bx;
        8'b1011_1101: vertical = 1'bx;
        8'b1011_1110: vertical = 1'bx;
        8'b1011_1111: vertical = 1'bx;

        8'b1100_0000: vertical = 1'bx;
        8'b1100_0001: vertical = 1'bx;
        8'b1100_0010: vertical = 1'bx;
        8'b1100_0011: vertical = 1'bx;
        8'b1100_0100: vertical = 1'bx;
        8'b1100_0101: vertical = 1'bx;
        8'b1100_0110: vertical = 1'bx;
        8'b1100_0111: vertical = 1'bx;
        8'b1100_1000: vertical = 1'bx;
        8'b1100_1001: vertical = 1'bx;
        8'b1100_1010: vertical = 1'bx;
        8'b1100_1011: vertical = 1'bx;
        8'b1100_1100: vertical = 1'bx;
        8'b1100_1101: vertical = 1'bx;
        8'b1100_1110: vertical = 1'bx;
        8'b1100_1111: vertical = 1'bx;

        8'b1101_0000: vertical = 1'bx;
        8'b1101_0001: vertical = 1'bx;
        8'b1101_0010: vertical = 1'bx;
        8'b1101_0011: vertical = 1'bx;
        8'b1101_0100: vertical = 1'bx;
        8'b1101_0101: vertical = 1'bx;
        8'b1101_0110: vertical = 1'bx;
        8'b1101_0111: vertical = 1'bx;
        8'b1101_1000: vertical = 1'bx;
        8'b1101_1001: vertical = 1'bx;
        8'b1101_1010: vertical = 1'bx;
        8'b1101_1011: vertical = 1'bx;
        8'b1101_1100: vertical = 1'bx;
        8'b1101_1101: vertical = 1'bx;
        8'b1101_1110: vertical = 1'bx;
        8'b1101_1111: vertical = 1'bx;

        8'b1110_0000: vertical = 1'bx;
        8'b1110_0001: vertical = 1'bx;
        8'b1110_0010: vertical = 1'bx;
        8'b1110_0011: vertical = 1'bx;
        8'b1110_0100: vertical = 1'bx;
        8'b1110_0101: vertical = 1'bx;
        8'b1110_0110: vertical = 1'bx;
        8'b1110_0111: vertical = 1'bx;
        8'b1110_1000: vertical = 1'bx;
        8'b1110_1001: vertical = 1'bx;
        8'b1110_1010: vertical = 1'bx;
        8'b1110_1011: vertical = 1'bx;
        8'b1110_1100: vertical = 1'bx;
        8'b1110_1101: vertical = 1'bx;
        8'b1110_1110: vertical = 1'bx;
        8'b1110_1111: vertical = 1'bx;

        8'b1111_0000: vertical = 1'bx;
        8'b1111_0001: vertical = 1'bx;
        8'b1111_0010: vertical = 1'bx;
        8'b1111_0011: vertical = 1'bx;
        8'b1111_0100: vertical = 1'bx;
        8'b1111_0101: vertical = 1'bx;
        8'b1111_0110: vertical = 1'bx;
        8'b1111_0111: vertical = 1'bx;
        8'b1111_1000: vertical = 1'bx;
        8'b1111_1001: vertical = 1'bx;
        8'b1111_1010: vertical = 1'bx;
        8'b1111_1011: vertical = 1'bx;
        8'b1111_1100: vertical = 1'bx;
        8'b1111_1101: vertical = 1'bx;
        8'b1111_1110: vertical = 1'bx;
        8'b1111_1111: vertical = 1'bx;

    endcase
end

endmodule
